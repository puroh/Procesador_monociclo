`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.10.2017 19:53:13
// Design Name: 
// Module Name: control_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module control_tb(
    input intruccion,
    output RegDest,
    output SaltoCond,
    output LeerMem,
    output MenmaReg,
    output ALUOp,
    output EscrMem,
    output FuenteALU,
    output escrReg
    );
endmodule
